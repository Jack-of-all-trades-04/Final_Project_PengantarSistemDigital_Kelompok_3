library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity wallet is
  port (
  );
end entity;

architecture rtl of wallet is

end architecture;
