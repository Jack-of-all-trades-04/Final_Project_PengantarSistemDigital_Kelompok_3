library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity block_header is
  port (
  );
end entity;

architecture rtl of block_header is

end architecture;
