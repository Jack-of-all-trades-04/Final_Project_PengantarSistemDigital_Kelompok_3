library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity hash64 is
  port (
  );
end entity;

architecture rtl of hash64 is

end architecture;
