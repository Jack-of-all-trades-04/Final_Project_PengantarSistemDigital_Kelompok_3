library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity top is
  port (
  );
end entity;

architecture rtl of top is

end architecture;
