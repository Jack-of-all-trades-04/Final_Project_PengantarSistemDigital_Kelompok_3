library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity miner is
  port (
  );
end entity;

architecture rtl of miner is

end architecture;
