library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity consensus_controller is
  port (
  );
end entity;

architecture rtl of consensus_controller is

end architecture;
